// start_cloud_hps_system.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module start_cloud_hps_system (
		input  wire        clk_clk,                       //      clk.clk
		input  wire [20:0] hex0_2_export,                 //   hex0_2.export
		input  wire [20:0] hex3_5_export,                 //   hex3_5.export
		inout  wire        hps_io_0_hps_io_sdio_inst_CMD, // hps_io_0.hps_io_sdio_inst_CMD
		inout  wire        hps_io_0_hps_io_sdio_inst_D0,  //         .hps_io_sdio_inst_D0
		inout  wire        hps_io_0_hps_io_sdio_inst_D1,  //         .hps_io_sdio_inst_D1
		output wire        hps_io_0_hps_io_sdio_inst_CLK, //         .hps_io_sdio_inst_CLK
		inout  wire        hps_io_0_hps_io_sdio_inst_D2,  //         .hps_io_sdio_inst_D2
		inout  wire        hps_io_0_hps_io_sdio_inst_D3,  //         .hps_io_sdio_inst_D3
		input  wire        hps_io_0_hps_io_uart0_inst_RX, //         .hps_io_uart0_inst_RX
		output wire        hps_io_0_hps_io_uart0_inst_TX, //         .hps_io_uart0_inst_TX
		output wire [3:0]  key_export,                    //      key.export
		input  wire [9:0]  ledr_export,                   //     ledr.export
		output wire [12:0] memory_mem_a,                  //   memory.mem_a
		output wire [2:0]  memory_mem_ba,                 //         .mem_ba
		output wire        memory_mem_ck,                 //         .mem_ck
		output wire        memory_mem_ck_n,               //         .mem_ck_n
		output wire        memory_mem_cke,                //         .mem_cke
		output wire        memory_mem_cs_n,               //         .mem_cs_n
		output wire        memory_mem_ras_n,              //         .mem_ras_n
		output wire        memory_mem_cas_n,              //         .mem_cas_n
		output wire        memory_mem_we_n,               //         .mem_we_n
		output wire        memory_mem_reset_n,            //         .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                 //         .mem_dq
		inout  wire        memory_mem_dqs,                //         .mem_dqs
		inout  wire        memory_mem_dqs_n,              //         .mem_dqs_n
		output wire        memory_mem_odt,                //         .mem_odt
		output wire        memory_mem_dm,                 //         .mem_dm
		input  wire        memory_oct_rzqin,              //         .oct_rzqin
		input  wire        reset_reset_n,                 //    reset.reset_n
		output wire [9:0]  sw_export                      //       sw.export
	);

	wire   [1:0] start_cloud_hps_h2f_lw_axi_master_awburst; // start_cloud_hps:h2f_lw_AWBURST -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awburst
	wire   [3:0] start_cloud_hps_h2f_lw_axi_master_arlen;   // start_cloud_hps:h2f_lw_ARLEN -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arlen
	wire   [3:0] start_cloud_hps_h2f_lw_axi_master_wstrb;   // start_cloud_hps:h2f_lw_WSTRB -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_wstrb
	wire         start_cloud_hps_h2f_lw_axi_master_wready;  // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_wready -> start_cloud_hps:h2f_lw_WREADY
	wire  [11:0] start_cloud_hps_h2f_lw_axi_master_rid;     // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_rid -> start_cloud_hps:h2f_lw_RID
	wire         start_cloud_hps_h2f_lw_axi_master_rready;  // start_cloud_hps:h2f_lw_RREADY -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_rready
	wire   [3:0] start_cloud_hps_h2f_lw_axi_master_awlen;   // start_cloud_hps:h2f_lw_AWLEN -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awlen
	wire  [11:0] start_cloud_hps_h2f_lw_axi_master_wid;     // start_cloud_hps:h2f_lw_WID -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_wid
	wire   [3:0] start_cloud_hps_h2f_lw_axi_master_arcache; // start_cloud_hps:h2f_lw_ARCACHE -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arcache
	wire         start_cloud_hps_h2f_lw_axi_master_wvalid;  // start_cloud_hps:h2f_lw_WVALID -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_wvalid
	wire  [20:0] start_cloud_hps_h2f_lw_axi_master_araddr;  // start_cloud_hps:h2f_lw_ARADDR -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_araddr
	wire   [2:0] start_cloud_hps_h2f_lw_axi_master_arprot;  // start_cloud_hps:h2f_lw_ARPROT -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arprot
	wire   [2:0] start_cloud_hps_h2f_lw_axi_master_awprot;  // start_cloud_hps:h2f_lw_AWPROT -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awprot
	wire  [31:0] start_cloud_hps_h2f_lw_axi_master_wdata;   // start_cloud_hps:h2f_lw_WDATA -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_wdata
	wire         start_cloud_hps_h2f_lw_axi_master_arvalid; // start_cloud_hps:h2f_lw_ARVALID -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arvalid
	wire   [3:0] start_cloud_hps_h2f_lw_axi_master_awcache; // start_cloud_hps:h2f_lw_AWCACHE -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awcache
	wire  [11:0] start_cloud_hps_h2f_lw_axi_master_arid;    // start_cloud_hps:h2f_lw_ARID -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arid
	wire   [1:0] start_cloud_hps_h2f_lw_axi_master_arlock;  // start_cloud_hps:h2f_lw_ARLOCK -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arlock
	wire   [1:0] start_cloud_hps_h2f_lw_axi_master_awlock;  // start_cloud_hps:h2f_lw_AWLOCK -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awlock
	wire  [20:0] start_cloud_hps_h2f_lw_axi_master_awaddr;  // start_cloud_hps:h2f_lw_AWADDR -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awaddr
	wire   [1:0] start_cloud_hps_h2f_lw_axi_master_bresp;   // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_bresp -> start_cloud_hps:h2f_lw_BRESP
	wire         start_cloud_hps_h2f_lw_axi_master_arready; // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arready -> start_cloud_hps:h2f_lw_ARREADY
	wire  [31:0] start_cloud_hps_h2f_lw_axi_master_rdata;   // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_rdata -> start_cloud_hps:h2f_lw_RDATA
	wire         start_cloud_hps_h2f_lw_axi_master_awready; // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awready -> start_cloud_hps:h2f_lw_AWREADY
	wire   [1:0] start_cloud_hps_h2f_lw_axi_master_arburst; // start_cloud_hps:h2f_lw_ARBURST -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arburst
	wire   [2:0] start_cloud_hps_h2f_lw_axi_master_arsize;  // start_cloud_hps:h2f_lw_ARSIZE -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_arsize
	wire         start_cloud_hps_h2f_lw_axi_master_bready;  // start_cloud_hps:h2f_lw_BREADY -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_bready
	wire         start_cloud_hps_h2f_lw_axi_master_rlast;   // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_rlast -> start_cloud_hps:h2f_lw_RLAST
	wire         start_cloud_hps_h2f_lw_axi_master_wlast;   // start_cloud_hps:h2f_lw_WLAST -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_wlast
	wire   [1:0] start_cloud_hps_h2f_lw_axi_master_rresp;   // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_rresp -> start_cloud_hps:h2f_lw_RRESP
	wire  [11:0] start_cloud_hps_h2f_lw_axi_master_awid;    // start_cloud_hps:h2f_lw_AWID -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awid
	wire  [11:0] start_cloud_hps_h2f_lw_axi_master_bid;     // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_bid -> start_cloud_hps:h2f_lw_BID
	wire         start_cloud_hps_h2f_lw_axi_master_bvalid;  // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_bvalid -> start_cloud_hps:h2f_lw_BVALID
	wire   [2:0] start_cloud_hps_h2f_lw_axi_master_awsize;  // start_cloud_hps:h2f_lw_AWSIZE -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awsize
	wire         start_cloud_hps_h2f_lw_axi_master_awvalid; // start_cloud_hps:h2f_lw_AWVALID -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_awvalid
	wire         start_cloud_hps_h2f_lw_axi_master_rvalid;  // mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_rvalid -> start_cloud_hps:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_ledr_pio_s1_readdata;    // ledr_pio:readdata -> mm_interconnect_0:ledr_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_pio_s1_address;     // mm_interconnect_0:ledr_pio_s1_address -> ledr_pio:address
	wire         mm_interconnect_0_sw_pio_s1_chipselect;    // mm_interconnect_0:sw_pio_s1_chipselect -> sw_pio:chipselect
	wire  [31:0] mm_interconnect_0_sw_pio_s1_readdata;      // sw_pio:readdata -> mm_interconnect_0:sw_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_pio_s1_address;       // mm_interconnect_0:sw_pio_s1_address -> sw_pio:address
	wire         mm_interconnect_0_sw_pio_s1_write;         // mm_interconnect_0:sw_pio_s1_write -> sw_pio:write_n
	wire  [31:0] mm_interconnect_0_sw_pio_s1_writedata;     // mm_interconnect_0:sw_pio_s1_writedata -> sw_pio:writedata
	wire         mm_interconnect_0_key_pio_s1_chipselect;   // mm_interconnect_0:key_pio_s1_chipselect -> key_pio:chipselect
	wire  [31:0] mm_interconnect_0_key_pio_s1_readdata;     // key_pio:readdata -> mm_interconnect_0:key_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_key_pio_s1_address;      // mm_interconnect_0:key_pio_s1_address -> key_pio:address
	wire         mm_interconnect_0_key_pio_s1_write;        // mm_interconnect_0:key_pio_s1_write -> key_pio:write_n
	wire  [31:0] mm_interconnect_0_key_pio_s1_writedata;    // mm_interconnect_0:key_pio_s1_writedata -> key_pio:writedata
	wire  [31:0] mm_interconnect_0_hex0_2_pio_s1_readdata;  // HEX0_2_pio:readdata -> mm_interconnect_0:HEX0_2_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_2_pio_s1_address;   // mm_interconnect_0:HEX0_2_pio_s1_address -> HEX0_2_pio:address
	wire  [31:0] mm_interconnect_0_hex3_5_pio_s1_readdata;  // HEX3_5_pio:readdata -> mm_interconnect_0:HEX3_5_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_5_pio_s1_address;   // mm_interconnect_0:HEX3_5_pio_s1_address -> HEX3_5_pio:address
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [HEX0_2_pio:reset_n, HEX3_5_pio:reset_n, key_pio:reset_n, ledr_pio:reset_n, mm_interconnect_0:ledr_pio_reset_reset_bridge_in_reset_reset, sw_pio:reset_n]
	wire         rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> mm_interconnect_0:start_cloud_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         start_cloud_hps_h2f_reset_reset;           // start_cloud_hps:h2f_rst_n -> rst_controller_001:reset_in0

	start_cloud_hps_system_HEX0_2_pio hex0_2_pio (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_hex0_2_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hex0_2_pio_s1_readdata), //                    .readdata
		.in_port  (hex0_2_export)                             // external_connection.export
	);

	start_cloud_hps_system_HEX0_2_pio hex3_5_pio (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_hex3_5_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_hex3_5_pio_s1_readdata), //                    .readdata
		.in_port  (hex3_5_export)                             // external_connection.export
	);

	start_cloud_hps_system_key_pio key_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_key_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_pio_s1_readdata),   //                    .readdata
		.out_port   (key_export)                               // external_connection.export
	);

	start_cloud_hps_system_ledr_pio ledr_pio (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_ledr_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ledr_pio_s1_readdata), //                    .readdata
		.in_port  (ledr_export)                             // external_connection.export
	);

	start_cloud_hps_system_start_cloud_hps #(
		.F2S_Width (0),
		.S2F_Width (0)
	) start_cloud_hps (
		.mem_a                (memory_mem_a),                              //            memory.mem_a
		.mem_ba               (memory_mem_ba),                             //                  .mem_ba
		.mem_ck               (memory_mem_ck),                             //                  .mem_ck
		.mem_ck_n             (memory_mem_ck_n),                           //                  .mem_ck_n
		.mem_cke              (memory_mem_cke),                            //                  .mem_cke
		.mem_cs_n             (memory_mem_cs_n),                           //                  .mem_cs_n
		.mem_ras_n            (memory_mem_ras_n),                          //                  .mem_ras_n
		.mem_cas_n            (memory_mem_cas_n),                          //                  .mem_cas_n
		.mem_we_n             (memory_mem_we_n),                           //                  .mem_we_n
		.mem_reset_n          (memory_mem_reset_n),                        //                  .mem_reset_n
		.mem_dq               (memory_mem_dq),                             //                  .mem_dq
		.mem_dqs              (memory_mem_dqs),                            //                  .mem_dqs
		.mem_dqs_n            (memory_mem_dqs_n),                          //                  .mem_dqs_n
		.mem_odt              (memory_mem_odt),                            //                  .mem_odt
		.mem_dm               (memory_mem_dm),                             //                  .mem_dm
		.oct_rzqin            (memory_oct_rzqin),                          //                  .oct_rzqin
		.hps_io_sdio_inst_CMD (hps_io_0_hps_io_sdio_inst_CMD),             //            hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0  (hps_io_0_hps_io_sdio_inst_D0),              //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1  (hps_io_0_hps_io_sdio_inst_D1),              //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK (hps_io_0_hps_io_sdio_inst_CLK),             //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2  (hps_io_0_hps_io_sdio_inst_D2),              //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3  (hps_io_0_hps_io_sdio_inst_D3),              //                  .hps_io_sdio_inst_D3
		.hps_io_uart0_inst_RX (hps_io_0_hps_io_uart0_inst_RX),             //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX (hps_io_0_hps_io_uart0_inst_TX),             //                  .hps_io_uart0_inst_TX
		.h2f_rst_n            (start_cloud_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_lw_axi_clk       (clk_clk),                                   //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID          (start_cloud_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR        (start_cloud_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN         (start_cloud_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE        (start_cloud_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST       (start_cloud_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK        (start_cloud_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE       (start_cloud_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT        (start_cloud_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID       (start_cloud_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY       (start_cloud_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID           (start_cloud_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA         (start_cloud_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB         (start_cloud_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST         (start_cloud_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID        (start_cloud_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY        (start_cloud_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID           (start_cloud_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP         (start_cloud_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID        (start_cloud_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY        (start_cloud_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID          (start_cloud_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR        (start_cloud_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN         (start_cloud_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE        (start_cloud_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST       (start_cloud_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK        (start_cloud_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE       (start_cloud_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT        (start_cloud_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID       (start_cloud_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY       (start_cloud_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID           (start_cloud_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA         (start_cloud_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP         (start_cloud_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST         (start_cloud_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID        (start_cloud_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY        (start_cloud_hps_h2f_lw_axi_master_rready)   //                  .rready
	);

	start_cloud_hps_system_sw_pio sw_pio (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_sw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_pio_s1_readdata),   //                    .readdata
		.out_port   (sw_export)                               // external_connection.export
	);

	start_cloud_hps_system_mm_interconnect_0 mm_interconnect_0 (
		.start_cloud_hps_h2f_lw_axi_master_awid                                        (start_cloud_hps_h2f_lw_axi_master_awid),    //                                       start_cloud_hps_h2f_lw_axi_master.awid
		.start_cloud_hps_h2f_lw_axi_master_awaddr                                      (start_cloud_hps_h2f_lw_axi_master_awaddr),  //                                                                        .awaddr
		.start_cloud_hps_h2f_lw_axi_master_awlen                                       (start_cloud_hps_h2f_lw_axi_master_awlen),   //                                                                        .awlen
		.start_cloud_hps_h2f_lw_axi_master_awsize                                      (start_cloud_hps_h2f_lw_axi_master_awsize),  //                                                                        .awsize
		.start_cloud_hps_h2f_lw_axi_master_awburst                                     (start_cloud_hps_h2f_lw_axi_master_awburst), //                                                                        .awburst
		.start_cloud_hps_h2f_lw_axi_master_awlock                                      (start_cloud_hps_h2f_lw_axi_master_awlock),  //                                                                        .awlock
		.start_cloud_hps_h2f_lw_axi_master_awcache                                     (start_cloud_hps_h2f_lw_axi_master_awcache), //                                                                        .awcache
		.start_cloud_hps_h2f_lw_axi_master_awprot                                      (start_cloud_hps_h2f_lw_axi_master_awprot),  //                                                                        .awprot
		.start_cloud_hps_h2f_lw_axi_master_awvalid                                     (start_cloud_hps_h2f_lw_axi_master_awvalid), //                                                                        .awvalid
		.start_cloud_hps_h2f_lw_axi_master_awready                                     (start_cloud_hps_h2f_lw_axi_master_awready), //                                                                        .awready
		.start_cloud_hps_h2f_lw_axi_master_wid                                         (start_cloud_hps_h2f_lw_axi_master_wid),     //                                                                        .wid
		.start_cloud_hps_h2f_lw_axi_master_wdata                                       (start_cloud_hps_h2f_lw_axi_master_wdata),   //                                                                        .wdata
		.start_cloud_hps_h2f_lw_axi_master_wstrb                                       (start_cloud_hps_h2f_lw_axi_master_wstrb),   //                                                                        .wstrb
		.start_cloud_hps_h2f_lw_axi_master_wlast                                       (start_cloud_hps_h2f_lw_axi_master_wlast),   //                                                                        .wlast
		.start_cloud_hps_h2f_lw_axi_master_wvalid                                      (start_cloud_hps_h2f_lw_axi_master_wvalid),  //                                                                        .wvalid
		.start_cloud_hps_h2f_lw_axi_master_wready                                      (start_cloud_hps_h2f_lw_axi_master_wready),  //                                                                        .wready
		.start_cloud_hps_h2f_lw_axi_master_bid                                         (start_cloud_hps_h2f_lw_axi_master_bid),     //                                                                        .bid
		.start_cloud_hps_h2f_lw_axi_master_bresp                                       (start_cloud_hps_h2f_lw_axi_master_bresp),   //                                                                        .bresp
		.start_cloud_hps_h2f_lw_axi_master_bvalid                                      (start_cloud_hps_h2f_lw_axi_master_bvalid),  //                                                                        .bvalid
		.start_cloud_hps_h2f_lw_axi_master_bready                                      (start_cloud_hps_h2f_lw_axi_master_bready),  //                                                                        .bready
		.start_cloud_hps_h2f_lw_axi_master_arid                                        (start_cloud_hps_h2f_lw_axi_master_arid),    //                                                                        .arid
		.start_cloud_hps_h2f_lw_axi_master_araddr                                      (start_cloud_hps_h2f_lw_axi_master_araddr),  //                                                                        .araddr
		.start_cloud_hps_h2f_lw_axi_master_arlen                                       (start_cloud_hps_h2f_lw_axi_master_arlen),   //                                                                        .arlen
		.start_cloud_hps_h2f_lw_axi_master_arsize                                      (start_cloud_hps_h2f_lw_axi_master_arsize),  //                                                                        .arsize
		.start_cloud_hps_h2f_lw_axi_master_arburst                                     (start_cloud_hps_h2f_lw_axi_master_arburst), //                                                                        .arburst
		.start_cloud_hps_h2f_lw_axi_master_arlock                                      (start_cloud_hps_h2f_lw_axi_master_arlock),  //                                                                        .arlock
		.start_cloud_hps_h2f_lw_axi_master_arcache                                     (start_cloud_hps_h2f_lw_axi_master_arcache), //                                                                        .arcache
		.start_cloud_hps_h2f_lw_axi_master_arprot                                      (start_cloud_hps_h2f_lw_axi_master_arprot),  //                                                                        .arprot
		.start_cloud_hps_h2f_lw_axi_master_arvalid                                     (start_cloud_hps_h2f_lw_axi_master_arvalid), //                                                                        .arvalid
		.start_cloud_hps_h2f_lw_axi_master_arready                                     (start_cloud_hps_h2f_lw_axi_master_arready), //                                                                        .arready
		.start_cloud_hps_h2f_lw_axi_master_rid                                         (start_cloud_hps_h2f_lw_axi_master_rid),     //                                                                        .rid
		.start_cloud_hps_h2f_lw_axi_master_rdata                                       (start_cloud_hps_h2f_lw_axi_master_rdata),   //                                                                        .rdata
		.start_cloud_hps_h2f_lw_axi_master_rresp                                       (start_cloud_hps_h2f_lw_axi_master_rresp),   //                                                                        .rresp
		.start_cloud_hps_h2f_lw_axi_master_rlast                                       (start_cloud_hps_h2f_lw_axi_master_rlast),   //                                                                        .rlast
		.start_cloud_hps_h2f_lw_axi_master_rvalid                                      (start_cloud_hps_h2f_lw_axi_master_rvalid),  //                                                                        .rvalid
		.start_cloud_hps_h2f_lw_axi_master_rready                                      (start_cloud_hps_h2f_lw_axi_master_rready),  //                                                                        .rready
		.clk_0_clk_clk                                                                 (clk_clk),                                   //                                                               clk_0_clk.clk
		.ledr_pio_reset_reset_bridge_in_reset_reset                                    (rst_controller_reset_out_reset),            //                                    ledr_pio_reset_reset_bridge_in_reset.reset
		.start_cloud_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),        // start_cloud_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.HEX0_2_pio_s1_address                                                         (mm_interconnect_0_hex0_2_pio_s1_address),   //                                                           HEX0_2_pio_s1.address
		.HEX0_2_pio_s1_readdata                                                        (mm_interconnect_0_hex0_2_pio_s1_readdata),  //                                                                        .readdata
		.HEX3_5_pio_s1_address                                                         (mm_interconnect_0_hex3_5_pio_s1_address),   //                                                           HEX3_5_pio_s1.address
		.HEX3_5_pio_s1_readdata                                                        (mm_interconnect_0_hex3_5_pio_s1_readdata),  //                                                                        .readdata
		.key_pio_s1_address                                                            (mm_interconnect_0_key_pio_s1_address),      //                                                              key_pio_s1.address
		.key_pio_s1_write                                                              (mm_interconnect_0_key_pio_s1_write),        //                                                                        .write
		.key_pio_s1_readdata                                                           (mm_interconnect_0_key_pio_s1_readdata),     //                                                                        .readdata
		.key_pio_s1_writedata                                                          (mm_interconnect_0_key_pio_s1_writedata),    //                                                                        .writedata
		.key_pio_s1_chipselect                                                         (mm_interconnect_0_key_pio_s1_chipselect),   //                                                                        .chipselect
		.ledr_pio_s1_address                                                           (mm_interconnect_0_ledr_pio_s1_address),     //                                                             ledr_pio_s1.address
		.ledr_pio_s1_readdata                                                          (mm_interconnect_0_ledr_pio_s1_readdata),    //                                                                        .readdata
		.sw_pio_s1_address                                                             (mm_interconnect_0_sw_pio_s1_address),       //                                                               sw_pio_s1.address
		.sw_pio_s1_write                                                               (mm_interconnect_0_sw_pio_s1_write),         //                                                                        .write
		.sw_pio_s1_readdata                                                            (mm_interconnect_0_sw_pio_s1_readdata),      //                                                                        .readdata
		.sw_pio_s1_writedata                                                           (mm_interconnect_0_sw_pio_s1_writedata),     //                                                                        .writedata
		.sw_pio_s1_chipselect                                                          (mm_interconnect_0_sw_pio_s1_chipselect)     //                                                                        .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~start_cloud_hps_h2f_reset_reset),   // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
